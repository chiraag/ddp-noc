typedef 3 Degree;
typedef 7 TotalNodes;

Integer incidence[3] = {
  0, 1, 3
};



